module Serial_32bits_add_sub();
	
	output [31:0] result;
	output overflow, Cout;
	input  [31:0] in1, in2;
	input  [1:0] OP; 






endmodule