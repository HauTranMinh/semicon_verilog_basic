module count_down_underflow_pclk2();

	

endmodule
